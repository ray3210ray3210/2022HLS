defparam AESL_inst_example.proc_1_U0.data_channel1_U.DEPTH = 'd10;
defparam AESL_inst_example.proc_1_U0.data_channel1_U.ADDR_WIDTH = 'd4;
defparam AESL_inst_example.data_channel2_U.DEPTH = 'd1;
defparam AESL_inst_example.data_channel2_U.ADDR_WIDTH = 'd0;
defparam AESL_inst_example.proc_1_U0.data_channel2_U.DEPTH = 'd1;
defparam AESL_inst_example.proc_1_U0.data_channel2_U.ADDR_WIDTH = 'd0;
defparam AESL_inst_example.proc_2_U0.data_channel2_U.DEPTH = 'd1;
defparam AESL_inst_example.proc_2_U0.data_channel2_U.ADDR_WIDTH = 'd0;
